LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE WORK.EE_232_Q1.ALL;
USE WORK.EE_232_PACKG.ALL;
ENTITY ALU_4 IS
PORT ( A, B : IN STD_LOGIC_VECTOR(3 DOWNTO 0) ;
S : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
F : OUT STD_LOGIC_VECTOR(3 DOWNTO 0) ;
O : OUT STD_LOGIC);
END ALU_4;


ARCHITECTURE FUNC OF ALU_4 IS
SIGNAL Y0, Y1, Y2, Y3, Y4, Y5, Y6, Y8: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL Y7 : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL F0, F1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL O0, O1, O2 : STD_LOGIC;

BEGIN
-- AND OPERATIONS

U0 : AND_2 PORT MAP (A(0),B(0),Y0(0));
U1 : AND_2 PORT MAP (A(1),B(1),Y0(1));
U2 : AND_2 PORT MAP (A(2),B(2),Y0(2));
U3 : AND_2 PORT MAP (A(3),B(3),Y0(3));

-- OR OPERATIONS

U4 : OR_2 PORT MAP (A(0),B(0),Y1(0));
U5 : OR_2 PORT MAP (A(1),B(1),Y1(1));
U6 : OR_2 PORT MAP (A(2),B(2),Y1(2));
U7 : OR_2 PORT MAP (A(3),B(3),Y1(3));

-- NOT OPERATIONS

U8  : NOT_2 PORT MAP (A(0),Y2(0));
U9  : NOT_2 PORT MAP (A(1),Y2(1));
U10 : NOT_2 PORT MAP (A(2),Y2(2));
U11 : NOT_2 PORT MAP (A(3),Y2(3));

-- XOR OPERATIONS

U12 : XOR_2 PORT MAP (A(0),B(0),Y3(0));
U13 : XOR_2 PORT MAP (A(1),B(1),Y3(1));
U14 : XOR_2 PORT MAP (A(2),B(2),Y3(2));
U15 : XOR_2 PORT MAP (A(3),B(3),Y3(3));


-- ADDITION OPERATIONS

AO : SUB_4 PORT MAP (A(0), A(1), A(2), A(3), B(0), B(1), B(2), B(3), S(0), Y4(0), Y4(1), Y4(2), Y4(3), O0); 

-- SUBTRACTION OPERATION

A1 : SUB_4 PORT MAP (A(0), A(1), A(2), A(3), B(0), B(1), B(2), B(3), S(0), Y5(0), Y5(1), Y5(2), Y5(3), O1); 

-- SUBTRACTION OPERATION

A2 : SUB_4 PORT MAP (B(0), B(1), B(2), B(3), A(0), A(1), A(2), A(3), S(1), Y6(0), Y6(1), Y6(2), Y6(3), O2); 

-- MULTIPLIcation operations
A3 : MULTIPLY_4 PORT MAP (A, B, Y7(0), Y7(1), Y7(2), Y7(3), Y7(4), Y7(5), Y7(6), Y7(7));


Y8(0) <= Y7(0);
Y8(1) <= Y7(1);
Y8(2) <= Y7(2);
Y8(3) <= Y7(3);

--  UNIT CONTROL 1

MO : mux_16_4 PORT MAP (Y4, Y5, Y6, Y0, S(1 DOWNTO 0), F0);

--  UNIT CONTROL 2

M1 : mux_16_4 PORT MAP (Y1, Y3, Y2, Y8, S(1 DOWNTO 0), F1);

-- OVERALL UNIT CONTROL

M2 : mux_2_1 PORT MAP (F0(0), F1(0), S(2), F(0));
M3 : mux_2_1 PORT MAP (F0(1), F1(1), S(2), F(1));
M4 : mux_2_1 PORT MAP (F0(2), F1(2), S(2), F(2));
M5 : mux_2_1 PORT MAP (F0(3), F1(3), S(2), F(3));

-- OVERFLOW CONTROL

M6 : MUX_8_1 PORT MAP (O0, O1, O2, '0', '0', '0', '0', Y7(4), S, O);

END ARCHITECTURE;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY NOT_2 IS
	PORT (I0: IN STD_LOGIC;
			O0 : OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE FUNC OF NOT_2 IS
BEGIN
	O0 <= NOT I0;
END FUNC;
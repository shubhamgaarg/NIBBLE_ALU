library ieee;
use ieeE.std_logic_1164.all;
USE WORK.EE_232_Q1.ALL;
USE WORK.EE_232_PACKG.ALL;
entity SUB_4 is 
port (A0,A1,A2,A3,B0,B1,B2,B3,AS : IN std_logic;
S0,S1,S2,S3,CO :OUT STD_LOGIC);
END ENTITY;
ARCHITECTURE FUNC OF SUB_4 IS 
SIGNAL M0,M1,M2,M3 : STD_LOGIC;
BEGIN 
U0 : XOR_2 PORT MAP (B0,AS,M0);
U1 : XOR_2 PORT MAP (B1,AS,M1);
U2 : XOR_2 PORT MAP (B2,AS,M2);
U3 : XOR_2 PORT MAP (B3,AS,M3);

F0 : FOUR_BIT_ADDER PORT MAP (A0,A1,A2,A3,M0,M1,M2,M3,AS,S0,S1,S2,S3,CO);
END FUNC;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE WORK.EE_232_PACKG.ALL;
ENTITY MUX_8_1 IS 
PORT (X0, X1, X2, X3, X4, X5, X6, X7 : IN  STD_LOGIC;
      S : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		Y : OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE FUNC OF MUX_8_1 IS
SIGNAL A,B : STD_LOGIC;
BEGIN
M0 : MUX_4_1 PORT MAP (X0, X1, X2, X3, S(1 DOWNTO 0), A);
M1 : MUX_4_1 PORT MAP (X4, X5, X6, X7, S(1 DOWNTO 0), B);
M2 : MUX_2_1 PORT MAP (A, B, S(2), Y);
END ARCHITECTURE; 
